module FSM();

endmodule
