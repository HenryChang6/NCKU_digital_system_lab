module vga_pic(

);


endmodule